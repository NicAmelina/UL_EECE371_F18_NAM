module test123; 
	reg A, B; 
	wire cout, c, acc;
	CB awful(A, B, c, cout, acc);
	initial
		begin
			A = 8'b00000001; B = 8'b00000110; 
			#20 A = 8'b00000001; B = 8'b01100100;
			#20 A = 8'b00000001; B = 8'b01111111; 
			#20 A = 8'b00000101; B = 8'b00001010;
			#20 A = 8'b00000101; B = 8'b01100100;
			#20 A = 8'b00000101; B = 8'b01111111;
			#20 A = 8'b01100100; B = 8'b01100100;
			#20 A = 8'b01100100; B = 8'b01111111;
			#20 A = 8'b01111111; B = 8'b01111111;

			#100 $finish;
		end
endmodule 

